module NOT(A_b, A);
    output A_b;
    input A;

    nand G1(A_b, A);

endmodule
