module AND16(O, I1, I2);
    output [15:0]O;
    input [15:0]I1, [15:0]I2;

    and G1(O, I1, I2);

endmodule
